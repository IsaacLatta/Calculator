----------------------------------------------------------------------------------
-- Company: Digilent Inc 2011
-- Engineer: Michelle Yu  
-- Create Date:    17:05:39 08/23/2011 
--
-- Module Name:    PmodKYPD - Behavioral 
-- Project Name:  PmodKYPD
-- Target Devices: Nexys3
-- Tool versions: Xilinx ISE 13.2 
-- Description: 
--	This file defines a project that outputs the key pressed on the PmodKYPD to the seven segment display
--
-- Revision: 
-- Revision 0.01 - File Created
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;
--use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity PmodKYPD is
    Port ( 
			  clk : in  STD_LOGIC;
			  JA : inout  STD_LOGIC_VECTOR (7 downto 0); -- PmodKYPD is designed to be connected to JA
           an : out  STD_LOGIC_VECTOR (3 downto 0);   -- Controls which position of the seven segment display to display
           seg : out  STD_LOGIC_VECTOR (6 downto 0); -- digit to display on the seven segment display 
           led : out STD_LOGIC_VECTOR(3 downto 0);
           input_debug: out STD_LOGIC_VECTOR(3 downto 0));
end PmodKYPD;

architecture Behavioral of PmodKYPD is

component Decoder is
	Port (
			 clk : in  STD_LOGIC;
            Row : in  STD_LOGIC_VECTOR (3 downto 0);
			 Col : out  STD_LOGIC_VECTOR (3 downto 0);
          DecodeOut : out  STD_LOGIC_VECTOR (3 downto 0));
	end component;

component DisplayController is
    Port ( 
        clk : in STD_LOGIC;                       -- Clock signal
        DispVal : in  STD_LOGIC_VECTOR (15 downto 0); -- 16-bit value to display
        anode : out std_logic_vector(3 downto 0); -- Anode control for four digits
        segOut : out  STD_LOGIC_VECTOR (6 downto 0)  -- Segment outputs
    );
end component;


component alu is
    Port (
        clk: in STD_LOGIC;
        done: out STD_LOGIC;
        ready: in STD_LOGIC;
        a : in  STD_LOGIC_VECTOR (15 downto 0);  -- Operand a (16 bits)
        b : in  STD_LOGIC_VECTOR (15 downto 0);  -- Operand b (16 bits)
        opcode : in STD_LOGIC_VECTOR (3 downto 0);  -- Operation selector
        result : out STD_LOGIC_VECTOR (31 downto 0)  -- Result (32 bits)
    );
end component;

component Debounce is
    Port ( 
        clk : in STD_LOGIC;
        input : in STD_LOGIC_VECTOR(3 downto 0);
        debounced : out STD_LOGIC_VECTOR(3 downto 0);
        input_changed : out STD_LOGIC
    );
    end component;

signal state: unsigned(3 downto 0) := to_unsigned(0, 4);
    signal enable: STD_LOGIC := '0'; 

    signal Decode: STD_LOGIC_VECTOR (3 downto 0) := "0000";
    signal Debounced_Decode: STD_LOGIC_VECTOR (3 downto 0) := "0000";
    signal Input_Changed: STD_LOGIC := '0';

   
    signal opcode: STD_LOGIC_VECTOR (3 downto 0) := "0000";
    signal operand_a: STD_LOGIC_VECTOR (15 downto 0) := (others => '0');
    signal operand_b: STD_LOGIC_VECTOR (15 downto 0) := (others => '0');
    signal result: STD_LOGIC_VECTOR (31 downto 0);  -- For multiplication results
    signal operand_a_ready: STD_LOGIC := '0';
    signal operand_b_ready: STD_LOGIC := '0';

    signal compute: STD_LOGIC := '0';
    signal completed: STD_LOGIC := '0';
    signal completed_last: STD_LOGIC := '0';  -- To detect rising edge of 'completed'
begin
    C0: Decoder port map (clk=>clk, Row =>JA(7 downto 4), Col=>JA(3 downto 0), DecodeOut=> Decode);
    C1: DisplayController port map (
    clk => clk,
    DispVal => result(15 downto 0),  -- Adjust based on result size
    anode => an,
    segOut => seg
    );

    C2: alu port map (
    clk => clk,  -- Pass the clock signal
    done => completed,
    ready => compute,
    a => operand_a,
    b => operand_b,
    opcode => opcode,
    result => result
    );

    C3: Debounce port map (
        clk => clk, 
        input => Decode, 
        debounced => Debounced_Decode,
        input_changed => Input_Changed
    );
    
    led <= STD_LOGIC_VECTOR(state);
    input_debug <= Debounced_Decode;
    --opcode <= "0000";  -- Always addition
-- Modify main_process
main_process: process(clk)
    variable digit_value: unsigned(3 downto 0);
begin
    if rising_edge(clk) then
        completed_last <= completed;  -- Update the previous 'completed' state
        case state is 
            when to_unsigned(0, 4) =>  -- Wait for first digit of operand A
                compute <= '0';
                operand_a <= (others => '0');
                operand_a_ready <= '0';
                if Input_Changed = '1' and Debounced_Decode /= "0000" then
                    digit_value := unsigned(Debounced_Decode);
                    operand_a <= std_logic_vector(resize(unsigned(operand_a) * 10 + unsigned(digit_value), 16));
                    state <= to_unsigned(1, 4);
                end if;
                
              
            when to_unsigned(1, 4) =>  -- Accumulate digits for operand A
                if Input_Changed = '1' then
                    if Debounced_Decode /= "1111" then  -- Assuming "1111" is 'Enter' or continue
                        digit_value := unsigned(Debounced_Decode);
                        operand_a <= std_logic_vector(resize(unsigned(operand_a) * 10 + unsigned(digit_value), 16));
                    else
                        operand_a_ready <= '1';
                        state <= to_unsigned(2, 4);
                    end if;
                end if;
                
            when to_unsigned(2, 4) =>  -- Wait for operator
                if Input_Changed = '1' and Debounced_Decode >= "1010" and Debounced_Decode <= "1101" then
                    opcode <= Debounced_Decode;
                    state <= to_unsigned(3, 4);
                end if;
                
            when to_unsigned(3, 4) =>  -- Wait for first digit of operand B
                operand_b <= (others => '0');
                operand_b_ready <= '0';
                if Input_Changed = '1' and Debounced_Decode /= "0000" then
                    digit_value := unsigned(Debounced_Decode);
                    operand_b <= std_logic_vector(resize(unsigned(operand_b) * 10 + unsigned(digit_value), 16));
                    state <= to_unsigned(4, 4);
                end if;
                
            when to_unsigned(4, 4) =>  -- Accumulate digits for operand B
                if Input_Changed = '1' then
                    if Debounced_Decode /= "1111" then  -- Assuming "1111" is 'Enter' or continue
                        digit_value := unsigned(Debounced_Decode);
                        operand_b <= std_logic_vector(resize(unsigned(operand_b) * 10 + unsigned(digit_value), 16));
                    else
                        operand_b_ready <= '1';
                        compute <= '1';  -- Start computation
                        state <= to_unsigned(5, 4);
                    end if;
                end if;
                
            when to_unsigned(5, 4) =>  -- Computation state
                if completed = '1' and completed_last = '0' then  -- Detect rising edge
                    compute <= '0';  -- Deassert compute after computation
                    state <= to_unsigned(6, 4);
                end if;
                
            when to_unsigned(6, 4) =>  -- Display result state
                -- Result is displayed; wait for user to reset
                if Input_Changed = '1' then
                    operand_a <= (others => '0');
                    operand_b <= (others => '0');
                    opcode <= (others => '0');
                    operand_a_ready <= '0';
                    operand_b_ready <= '0';
                    state <= to_unsigned(0, 4);
                end if;
                
            when others =>
                state <= to_unsigned(8, 4);  -- Invalid state for debugging
        end case;
    end if;
end process;

end Behavioral;
